library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

use work.records.all;


package pmemContent is

   constant pmemc : pmem_t := (
         ("01010" & "000" & "0000" & "0000" & "0000" & "0000" & "0001" & "0000"), -- BRA.wo #16
         ("00000" & "000" & "0000" & "0000" & "0000" & "0000" & "0000" & "0000"), -- NOP
         ("01001" & "000" & "0000" & "0000" & "0000" & "0000" & "0000" & "0001"), -- BRA.wofr R1
         ("00000" & "000" & "0000" & "0000" & "0000" & "0000" & "0000" & "0000"), -- NOP
         
         ("00110" & "01100" & "00001" & "0" & "0000" & "0000" & "0000" & "0010"), -- CMP.c
         ("10000" & "0000" & "000" & "0000" & "0000" & "0000" & "0000" & "1000"), -- BRZ.a #8
         ("00000" & "000" & "0000" & "0000" & "0000" & "0000" & "0000" & "0000"), -- NOP
         ("00000" & "000" & "0000" & "0000" & "0000" & "0000" & "0000" & "0000"), -- NOP
         
         
         ("10100" & "0000" & "000" & "0000" & "0000" & "0000" & "0000" & "1100"), -- BNZ.a #12
         ("00000" & "000" & "0000" & "0000" & "0000" & "0000" & "0000" & "0000"), -- NOP
         ("00000" & "000" & "0000" & "0000" & "0000" & "0000" & "0000" & "0000"), -- NOP
         ("00000" & "000" & "0000" & "0000" & "0000" & "0000" & "0000" & "0000"), -- NOP
         
         ("00110" & "00001" & "00001" & "0" & "0000" & "0000" & "0000" & "0001"), -- ADD R1 #1
         ("10100" & "0000" & "000" & "0000" & "0000" & "0000" & "0001" & "0000"), -- BNZ.a #32
         ("00000" & "000" & "0000" & "0000" & "0000" & "0000" & "0000" & "0000"), -- NOP
         ("01000" & "000" & "0000" & "0000" & "0000" & "0000" & "0000" & "0000"), -- BRA.a #0
         
         ("11101" & "00001" & "00" & "0000" & "0000" & "0000" & "0000" & "0010"), -- LOAD.c R1 #2
         ("00000" & "000" & "0000" & "0000" & "0000" & "0000" & "0000" & "0000"), -- NOP
         ("00000" & "000" & "0000" & "0000" & "0000" & "0000" & "0000" & "0000"), -- NOP
         ("01000" & "000" & "0000" & "0000" & "0000" & "0000" & "0000" & "0010"), -- BRA.a #2
         
         ("00000" & "000" & "0000" & "0000" & "0000" & "0000" & "0000" & "0000"), -- NOP
         ("00000" & "000" & "0000" & "0000" & "0000" & "0000" & "0000" & "0000"), -- NOP
         ("00000" & "000" & "0000" & "0000" & "0000" & "0000" & "0000" & "0000"), -- NOP
         ("00000" & "000" & "0000" & "0000" & "0000" & "0000" & "0000" & "0000"), -- NOP

      others =>
         ("00000" & "000" & "0000" & "0000" & "0000" & "0000" & "0000" & "0000")
      );
      
end pmemContent;
