library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

use work.Constants.all;

   --1 tile = 16x16 pixlar
   --30 tiles i x-led
   --17 tiles i y-led
   --30*17= tiles totalt på skärmen
   --dmem 16 bitar brett
   -- XXXX XXXX XXXX XXXX
   --Behöver 5 bitar för att peka ut rätt tile i tilemem
   -- Varje minnesplats i dmem får hålla reda på 3 tiles
   --1 vit
   --0 svart

package tilememContent is
   type tile_mem_c is array (0 to TILE_DIM - 1) of std_logic_vector(0 to TILE_DIM - 1);
   type tile_mem_t is array (0 to TILE_MEM_HEIGHT - 1) of tile_mem_c;

   constant tileMemoryContent : tile_mem_t := (
         --0
         (("0011111111111100"),
          ("0010000000001100"),
          ("0010000000010100"),
          ("0010000000100100"),
          ("0010000001000100"),
          ("0010000010000100"),
          ("0010000100000100"),
          ("0010001000000100"),
          ("0010010000000100"),
          ("0010100000000100"),
          ("0011000000000100"),
          ("0010000000000100"),
          ("0011111111111100"),
          ("0000000000000000"),
          ("0000000000000000"),
          ("0000000000000000")),
         --1
         (("0000000000000100"),
          ("0000000000000100"),
          ("0000000000000100"),
          ("0000000000000100"),
          ("0000000000000100"),
          ("0000000000000100"),
          ("0000000000000100"),
          ("0000000000000100"),
          ("0000000000000100"),
          ("0000000000000100"),
          ("0000000000000100"),
          ("0000000000000100"),
          ("0000000000000100"),
          ("0000000000000000"),
          ("0000000000000000"),
          ("0000000000000000")),
         --2
         (("0011111111111100"),
          ("0000000000000100"),
          ("0000000000000100"),
          ("0000000000000100"),
          ("0000000000000100"),
          ("0000000000000100"),
          ("0011111111111100"),
          ("0010000000000000"),
          ("0010000000000000"),
          ("0010000000000000"),
          ("0010000000000000"),
          ("0010000000000000"),
          ("0011111111111100"),
          ("0000000000000000"),
          ("0000000000000000"),
          ("0000000000000000")),
         --3
         (("0011111111111100"),
          ("0000000000000100"),
          ("0000000000000100"),
          ("0000000000000100"),
          ("0000000000000100"),
          ("0000000000000100"),
          ("0011111111111100"),
          ("0000000000000010"),
          ("0000000000000010"),
          ("0000000000000010"),
          ("0000000000000010"),
          ("0000000000000010"),
          ("0011111111111100"),
          ("0000000000000000"),
          ("0000000000000000"),
          ("0000000000000000")),
         --4
         (("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0011111111111100"),
          ("0000000000000100"),
          ("0000000000000100"),
          ("0000000000000100"),
          ("0000000000000100"),
          ("0000000000000100"),
          ("0000000000000100"),
          ("0000000000000000"),
          ("0000000000000000"),
          ("0000000000000000")),

         --5
         (("0011111111111100"),
          ("0010000000000000"),
          ("0010000000000000"),
          ("0010000000000000"),
          ("0010000000000000"),
          ("0010000000000000"),
          ("0011111111111100"),
          ("0000000000000100"),
          ("0000000000000100"),
          ("0000000000000100"),
          ("0000000000000100"),
          ("0000000000000100"),
          ("0011111111111100"),
          ("0000000000000000"),
          ("0000000000000000"),
          ("0000000000000000")),

         --6
         (("0011111111111100"),
          ("0010000000000000"),
          ("0010000000000000"),
          ("0010000000000000"),
          ("0010000000000000"),
          ("0010000000000000"),
          ("0011111111111100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0011111111111100"),
          ("0000000000000000"),
          ("0000000000000000"),
          ("0000000000000000")),

         --7
         (("0011111111111100"),
          ("0000000000000100"),
          ("0000000000000100"),
          ("0000000000000100"),
          ("0000000000000100"),
          ("0000000000000100"),
          ("0000000000000100"),
          ("0000000000000100"),
          ("0000000000000100"),
          ("0000000000000100"),
          ("0000000000000100"),
          ("0000000000000100"),
          ("0000000000000100"),
          ("0000000000000000"),
          ("0000000000000000"),
          ("0000000000000000")),

         --8
         (("0011111111111100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0011111111111100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0011111111111100"),
          ("0000000000000000"),
          ("0000000000000000"),
          ("0000000000000000")),

         --9
         (("0011111111111100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0011111111111100"),
          ("0000000000000100"),
          ("0000000000000100"),
          ("0000000000000100"),
          ("0000000000000100"),
          ("0000000000000100"),
          ("0000000000000100"),
          ("0000000000000000"),
          ("0000000000000000"),
          ("0000000000000000")),

         --A
         (("0001111111111000"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0011111111111100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0000000000000000"),
          ("0000000000000000"),
          ("0000000000000000")),

         --B
         (("0011111111110000"),
          ("0010000000001000"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000001000"),
          ("0011111111110000"),
          ("0010000000001000"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000001000"),
          ("0011111111110000"),
          ("0000000000000000"),
          ("0000000000000000"),
          ("0000000000000000")),

         --C
         (("0000111111111000"),
          ("0001000000000000"),
          ("0010000000000000"),
          ("0010000000000000"),
          ("0010000000000000"),
          ("0010000000000000"),
          ("0010000000000000"),
          ("0010000000000000"),
          ("0010000000000000"),
          ("0010000000000000"),
          ("0010000000000000"),
          ("0010000000000000"),
          ("0001111111111100"),
          ("0000000000000000"),
          ("0000000000000000"),
          ("0000000000000000")),

         --D
         (("0011111111110000"),
          ("0010000000001000"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000001000"),
          ("0011111111110000"),
          ("0000000000000000"),
          ("0000000000000000"),
          ("0000000000000000")),

         --E
         (("0011111111111100"),
          ("0010000000000000"),
          ("0010000000000000"),
          ("0010000000000000"),
          ("0010000000000000"),
          ("0010000000000000"),
          ("0011111111111100"),
          ("0010000000000000"),
          ("0010000000000000"),
          ("0010000000000000"),
          ("0010000000000000"),
          ("0010000000000000"),
          ("0011111111111100"),
          ("0000000000000000"),
          ("0000000000000000"),
          ("0000000000000000")),

         --F
         (("0011111111111100"),
          ("0010000000000000"),
          ("0010000000000000"),
          ("0010000000000000"),
          ("0010000000000000"),
          ("0010000000000000"),
          ("0011111111111100"),
          ("0010000000000000"),
          ("0010000000000000"),
          ("0010000000000000"),
          ("0010000000000000"),
          ("0010000000000000"),
          ("0010000000000000"),
          ("0000000000000000"),
          ("0000000000000000"),
          ("0000000000000000")),
         
         --H
         (("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0011111111111100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0000000000000000"),
          ("0000000000000000"),
          ("0000000000000000")),

         --I
         (("0000001110000000"),
          ("0000000100000000"),
          ("0000000100000000"),
          ("0000000100000000"),
          ("0000000100000000"),
          ("0000000100000000"),
          ("0000000100000000"),
          ("0000000100000000"),
          ("0000000100000000"),
          ("0000000100000000"),
          ("0000000100000000"),
          ("0000000100000000"),
          ("0000001110000000"),
          ("0000000000000000"),
          ("0000000000000000"),
          ("0000000000000000")),

         --I
         (("0010000000000000"),
          ("0010000000000000"),
          ("0010000000000000"),
          ("0010000000000000"),
          ("0010000000000000"),
          ("0010000000000000"),
          ("0010000000000000"),
          ("0010000000000000"),
          ("0010000000000000"),
          ("0010000000000000"),
          ("0010000000000000"),
          ("0010000000000000"),
          ("0011111111111100"),
          ("0000000000000000"),
          ("0000000000000000"),
          ("0000000000000000")),

         --N
         (("0010000000000100"),
          ("0011000000000100"),
          ("0010100000000100"),
          ("0010010000000100"),
          ("0010001000000100"),
          ("0010000100000100"),
          ("0010000100000100"),
          ("0010000010000100"),
          ("0010000001000100"),
          ("0010000000100100"),
          ("0010000000010100"),
          ("0010000000001100"),
          ("0010000000000100"),
          ("0000000000000000"),
          ("0000000000000000"),
          ("0000000000000000")),

         --O
         (("0000011111100000"),
          ("0000100000010000"),
          ("0001000000001000"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0001000000001000"),
          ("0000100000010000"),
          ("0000011111100000"),
          ("0000000000000000"),
          ("0000000000000000"),
          ("0000000000000000")),

         --P
         (("0011111111110000"),
          ("0010000000001000"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000001000"),
          ("0011111111110000"),
          ("0010000000000000"),
          ("0010000000000000"),
          ("0010000000000000"),
          ("0010000000000000"),
          ("0010000000000000"),
          ("0010000000000000"),
          ("0000000000000000"),
          ("0000000000000000"),
          ("0000000000000000")),

         --Q
         (("0000011111100000"),
          ("0000100000010000"),
          ("0001000000001000"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000100100"),
          ("0001000000011000"),
          ("0000100000011000"),
          ("0000011111100100"),
          ("0000000000000000"),
          ("0000000000000000"),
          ("0000000000000000")),

         --R
         (("0011111111110000"),
          ("0010000000001000"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000001000"),
          ("0011111111110000"),
          ("0010000000010000"),
          ("0010000000001000"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0000000000000000"),
          ("0000000000000000"),
          ("0000000000000000")),

         --S
         (("0000111111110000"),
          ("0001000000001000"),
          ("0010000000000100"),
          ("0010000000000000"),
          ("0001000000000000"),
          ("0000100000000000"),
          ("0000011111100000"),
          ("0000000000010000"),
          ("0000000000001000"),
          ("0000000000000100"),
          ("0010000000000100"),
          ("0001000000001000"),
          ("0000111111110000"),
          ("0000000000000000"),
          ("0000000000000000"),
          ("0000000000000000")),

         --T
         (("0011111111111100"),
          ("0000000100000000"),
          ("0000000100000000"),
          ("0000000100000000"),
          ("0000000100000000"),
          ("0000000100000000"),
          ("0000000100000000"),
          ("0000000100000000"),
          ("0000000100000000"),
          ("0000000100000000"),
          ("0000000100000000"),
          ("0000000100000000"),
          ("0000000100000000"),
          ("0000000000000000"),
          ("0000000000000000"),
          ("0000000000000000")),

         --U
         (("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0001000000001000"),
          ("0000100000010000"),
          ("0000011111100000"),
          ("0000000000000000"),
          ("0000000000000000"),
          ("0000000000000000")),

         --V
         (("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0001000000001000"),
          ("0000100000010000"),
          ("0000010000100000"),
          ("0000001001000000"),
          ("0000000110000000"),
          ("0000000000000000"),
          ("0000000000000000"),
          ("0000000000000000")),

         --w
         (("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0010000110000100"),
          ("0010000110000100"),
          ("0010000110000100"),
          ("0001000110001000"),
          ("0000101001010000"),
          ("0000010000100000"),
          ("0000000000000000"),
          ("0000000000000000"),
          ("0000000000000000")),

         --Y
         (("0010000000000100"),
          ("0010000000000100"),
          ("0010000000000100"),
          ("0001000000001000"),
          ("0000100000110000"),
          ("0000011111000000"),
          ("0000000100000000"),
          ("0000000100000000"),
          ("0000000100000000"),
          ("0000000100000000"),
          ("0000000100000000"),
          ("0000000100000000"),
          ("0000000100000000"),
          ("0000000100000000"),
          ("0000000000000000"),
          ("0000000000000000")),

         --space
         (("0000000000000000"),
          ("0000000000000000"),
          ("0000000000000000"),
          ("0000000000000000"),
          ("0000000000000000"),
          ("0000000000000000"),
          ("0000000000000000"),
          ("0000000000000000"),
          ("0000000000000000"),
          ("0000000000000000"),
          ("0000000000000000"),
          ("0000000000000000"),
          ("0000000000000000"),
          ("0000000000000000"),
          ("0000000000000000"),
          ("0000000000000000")),

         --colon :
         (("0000000000000000"),
          ("0001100000000000"),
          ("0001100000000000"),
          ("0000000000000000"),
          ("0000000000000000"),
          ("0000000000000000"),
          ("0001100000000000"),
          ("0001100000000000"),
          ("0000000000000000"),
          ("0000000000000000"),
          ("0000000000000000"),
          ("0000000000000000"),
          ("0000000000000000"),
          ("0000000000000000"),
          ("0000000000000000"),
          ("0000000000000000"))
      );
      
end tilememContent;
