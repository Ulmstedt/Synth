library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

use work.records.all;


package pmemContent is
   constant pmemc : pmem_t := (
         ("11000" & "00000" & "00" & "0000" & "0000" & "0000" & "0000" & "1110"),
         ("00000" & "000" & "0000" & "0000" & "0000" & "0000" & "0000" & "0000"),
         ("00000" & "000" & "0000" & "0000" & "0000" & "0000" & "0000" & "0000"),
         ("00000" & "000" & "0000" & "0000" & "0000" & "0000" & "0000" & "0000"),
         ("00000" & "000" & "0000" & "0000" & "0000" & "0000" & "0000" & "0000"),
         ("00000" & "000" & "0000" & "0000" & "0000" & "0000" & "0000" & "0000"),
         ("00000" & "000" & "0000" & "0000" & "0000" & "0000" & "0000" & "0000"),
         ("00000" & "000" & "0000" & "0000" & "0000" & "0000" & "0000" & "0000"),
      others =>
         ("00000" & "000" & "0000" & "0000" & "0000" & "0000" & "0000" & "0000")
      );
      
end pmemContent;