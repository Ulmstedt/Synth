library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

use work.records.all;
use work.Constants.all;


package memContent is
   constant memc : mem_t := (
      -- Wavetables (calculated in advance as: freq * wavetable_length / sample rate
      ("0000000010110000"), -- C0
      ("0000000010111010"),
      ("0000000011000101"),
      ("0000000011010001"),
      ("0000000011011101"),
      ("0000000011101010"),
      ("0000000011111000"),
      ("0000000100000111"),
      ("0000000100010111"),
      ("0000000100100111"),
      ("0000000100111001"),
      ("0000000101001011"),
      ("0000000101011111"),
      ("0000000101110100"),
      ("0000000110001010"),
      ("0000000110100010"),
      ("0000000110111010"),
      ("0000000111010101"),
      ("0000000111110000"),
      ("0000001000001110"),
      ("0000001000101101"),
      ("0000001001001111"),
      ("0000001001110010"),
      ("0000001010010111"),
      ("0000001010111110"),
      ("0000001011101000"),
      ("0000001100010100"),
      ("0000001101000011"),
      ("0000001101110101"),
      ("0000001110101010"),
      ("0000001111100001"),
      ("0000010000011100"),
      ("0000010001011011"),
      ("0000010010011101"),
      ("0000010011100100"),
      ("0000010100101110"),
      ("0000010101111100"),
      ("0000010111010000"),
      ("0000011000101000"),
      ("0000011010000111"),
      ("0000011011101010"),
      ("0000011101010011"),
      ("0000011111000010"),
      ("0000100000111001"),
      ("0000100010110110"),
      ("0000100100111010"),
      ("0000100111000111"),
      ("0000101001011100"),
      ("0000101011111001"),
      ("0000101110100000"),
      ("0000110001010001"),
      ("0000110100001101"),
      ("0000110111010011"),
      ("0000111010100110"),
      ("0000111110000100"),
      ("0001000001110001"),
      ("0001000101101100"),
      ("0001001001110100"),
      ("0001001110001110"),
      ("0001010010110111"),
      ("0001010111110010"),
      ("0001011100111111"),
      ("0001100010100001"),
      ("0001101000011011"),
      ("0001101110100110"),
      ("0001110101001101"),
      ("0001111100001000"),
      ("0010000011100010"),
      ("0010001011011000"),
      ("0010010011101001"),
      ("0010011100011100"),
      ("0010100101101111"),
      ("0010101111100100"),
      ("0010111001111110"),
      ("0011000101000010"),
      ("0011010000110110"),
      ("0011011101001100"),
      ("0011101010011010"),
      ("0011111000010000"),
      ("0100000111000100"),
      ("0100010110110000"),
      ("0100100111010010"),
      ("0100111000111001"),
      ("0101001011011110"), -- B6
      -- 64 step square wave
      ("1000000001000000"), 
      ("1000000001000000"), 
      ("1000000001000000"), 
      ("1000000001000000"), 
      ("1000000001000000"), 
      ("1000000001000000"), 
      ("1000000001000000"), 
      ("1000000001000000"), 
      ("1000000001000000"), 
      ("1000000001000000"), 
      ("1000000001000000"), 
      ("1000000001000000"), 
      ("1000000001000000"), 
      ("1000000001000000"), 
      ("1000000001000000"), 
      ("1000000001000000"), 
      ("1000000001000000"), 
      ("1000000001000000"), 
      ("1000000001000000"), 
      ("1000000001000000"), 
      ("1000000001000000"), 
      ("1000000001000000"), 
      ("1000000001000000"), 
      ("1000000001000000"), 
      ("1000000001000000"), 
      ("1000000001000000"), 
      ("1000000001000000"), 
      ("1000000001000000"), 
      ("1000000001000000"), 
      ("1000000001000000"), 
      ("1000000001000000"), 
      ("1000000001000000"), 
      ("0111111111000000"), 
      ("0111111111000000"), 
      ("0111111111000000"), 
      ("0111111111000000"), 
      ("0111111111000000"), 
      ("0111111111000000"), 
      ("0111111111000000"), 
      ("0111111111000000"), 
      ("0111111111000000"), 
      ("0111111111000000"), 
      ("0111111111000000"), 
      ("0111111111000000"), 
      ("0111111111000000"), 
      ("0111111111000000"), 
      ("0111111111000000"), 
      ("0111111111000000"), 
      ("0111111111000000"), 
      ("0111111111000000"), 
      ("0111111111000000"), 
      ("0111111111000000"), 
      ("0111111111000000"), 
      ("0111111111000000"), 
      ("0111111111000000"), 
      ("0111111111000000"), 
      ("0111111111000000"), 
      ("0111111111000000"), 
      ("0111111111000000"), 
      ("0111111111000000"), 
      ("0111111111000000"), 
      ("0111111111000000"), 
      ("0111111111000000"), 
      ("0111111111000000"), 
      -- 64 step sin wave
      ("0000110010000101"), 
      ("0001100011101100"), 
      ("0010010100010101"), 
      ("0011000011100011"), 
      ("0011110000111000"), 
      ("0100011011111001"), 
      ("0101000100001011"), 
      ("0101101001010101"), 
      ("0110001011000000"), 
      ("0110101000111000"), 
      ("0111000010101010"), 
      ("0111011000000110"), 
      ("0111101000111111"), 
      ("0111110101001011"), 
      ("0111111100100010"), 
      ("0111111111000000"), 
      ("0111111100100010"), 
      ("0111110101001011"), 
      ("0111101000111111"), 
      ("0111011000000110"), 
      ("0111000010101010"), 
      ("0110101000111000"), 
      ("0110001011000000"), 
      ("0101101001010101"), 
      ("0101000100001011"), 
      ("0100011011111001"), 
      ("0011110000111000"), 
      ("0011000011100011"), 
      ("0010010100010101"), 
      ("0001100011101100"), 
      ("0000110010000101"), 
      ("0000000000000000"), 
      ("1111001101111010"), 
      ("1110011100010011"), 
      ("1101101011101010"), 
      ("1100111100011100"), 
      ("1100001111000111"), 
      ("1011100100000110"), 
      ("1010111011110100"), 
      ("1010010110101010"), 
      ("1001110100111111"), 
      ("1001010111000111"), 
      ("1000111101010101"), 
      ("1000100111111001"), 
      ("1000010111000000"), 
      ("1000001010110100"), 
      ("1000000011011101"), 
      ("1000000001000000"), 
      ("1000000011011101"), 
      ("1000001010110100"), 
      ("1000010111000000"), 
      ("1000100111111001"), 
      ("1000111101010101"), 
      ("1001010111000111"), 
      ("1001110100111111"), 
      ("1010010110101010"), 
      ("1010111011110100"), 
      ("1011100100000110"), 
      ("1100001111000111"), 
      ("1100111100011100"), 
      ("1101101011101010"), 
      ("1110011100010011"), 
      ("1111001101111010"), 
      ("1111111111111111"), 
      -- 64 step saw wave
      ("0111101111000010"), 
      ("0111011111000100"), 
      ("0111001111000110"), 
      ("0110111111001000"), 
      ("0110101111001010"), 
      ("0110011111001100"), 
      ("0110001111001110"), 
      ("0101111111010000"), 
      ("0101101111010010"), 
      ("0101011111010100"), 
      ("0101001111010110"), 
      ("0100111111011000"), 
      ("0100101111011010"), 
      ("0100011111011100"), 
      ("0100001111011110"), 
      ("0011111111100000"), 
      ("0011101111100010"), 
      ("0011011111100100"), 
      ("0011001111100110"), 
      ("0010111111101000"), 
      ("0010101111101010"), 
      ("0010011111101100"), 
      ("0010001111101110"), 
      ("0001111111110000"), 
      ("0001101111110010"), 
      ("0001011111110100"), 
      ("0001001111110110"), 
      ("0000111111111000"), 
      ("0000101111111010"), 
      ("0000011111111100"), 
      ("0000001111111110"), 
      ("0000000000000000"), 
      ("1111110000000010"), 
      ("1111100000000100"), 
      ("1111010000000110"), 
      ("1111000000001000"), 
      ("1110110000001010"), 
      ("1110100000001100"), 
      ("1110010000001110"), 
      ("1110000000010000"), 
      ("1101110000010010"), 
      ("1101100000010100"), 
      ("1101010000010110"), 
      ("1101000000011000"), 
      ("1100110000011010"), 
      ("1100100000011100"), 
      ("1100010000011110"), 
      ("1100000000100000"), 
      ("1011110000100010"), 
      ("1011100000100100"), 
      ("1011010000100110"), 
      ("1011000000101000"), 
      ("1010110000101010"), 
      ("1010100000101100"), 
      ("1010010000101110"), 
      ("1010000000110000"), 
      ("1001110000110010"), 
      ("1001100000110100"), 
      ("1001010000110110"), 
      ("1001000000111000"), 
      ("1000110000111010"), 
      ("1000100000111100"), 
      ("1000010000111110"), 
      ("1000000001000000"),
      -- Cordic
      --TILE_MAP_OFFSET =>
      --   ("0000" & "0001" & "0000" & "0001" ),
      --TILE_MAP_OFFSET + 4 =>
      --   ("0000" & "0001" & "0000" & "0001" ),
      others =>
         ("0000" & "0000" & "0000" & "0000" )
      );
      
end memContent;
