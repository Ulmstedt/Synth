library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

use work.records.all;


package pmemContent is
   constant pmemc : pmem_t := (
         ("00000" & "00000" & "00" & "0000" & "0000" & "0000" & "0000" & "0000"),
         ("11100" & "000" & "0100" & "0000" & "0000" & "0000" & "0000" & "0000"),
         ("11100" & "000" & "1000" & "0000" & "0000" & "0000" & "0000" & "0001"),
         ("11100" & "000" & "1100" & "0000" & "0000" & "0000" & "0000" & "0010"),
         ("00000" & "000" & "0000" & "0000" & "0000" & "0000" & "0000" & "0000"),
         ("00000" & "000" & "0000" & "0000" & "0000" & "0000" & "0000" & "0000"),
      others =>
         ("00000" & "000" & "0000" & "0000" & "0000" & "0000" & "0000" & "0000")
      );
      
end pmemContent;
