library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

use work.records.all;


package pmemContent is

   constant pmemc : pmem_t := (

("11101100100000000000100000000000"),
("01000000000000000000000000001010"),
("00000000000000000000000000000000"),
("00000000000000000000000000000000"),
("00000000000000000000000000000000"),
("00000000000000000000000000000000"),
("10000010100000000000000000011101"),
("00000000000000000000000000000000"),
("01000000000000000000000000000001"),
("00000000000000000000000000000000"),
("10100011100000000000000000000011"),
("00000000000000000000000000000000"),
("00100000000000000000000000011101"),
("00110010000000000000000011111111"),
("00100000010000000000000000011110"),
("11101000100000000000001000000000"),
("00110011000000100000000000000000"),
("10000000000000000000000000011000"),
("00000000000000000000000000000000"),
("11011000000000000001000000000000"),
("11101001000000000000000000000001"),
("11011000000000010001000000000100"),
("01000000000000000000000000011011"),
("00000000000000000000000000000000"),
("11101001000000000000000000000000"),
("00000000000000000000000000000000"),
("11011000000000000001000000000100"),
("01000000000000000000000000000011"),
("00000000000000000000000000000000"),
("11101100100000000000100000000000"),
("11101000100000000000001000000000"),
("11111000000001000000000000000000"),
("00110011000000000000000000000000"),
("10000000000000000000000000101010"),
("11111001100000000000000000000000"),
("11111001110001000000000000000001"),
("00110000100011100000000000000001"),
("00101100010011000000000000000111"),
("00110000100001000000000000000001"),
("11011000000000000001000000000111"),
("00110010000011000000000000111111"),
("11111111110011000000000011010100"),
("01000000000000000000000000001000"),
("00000000000000000000000000000000"),

         -- Simple sound test
         --("11101111110000000000111111111111"),
         --("11101100100000001111110111101000"),
         --("10100010100000000000000000000010"),
         --("00000000000000000000000000000000"),
         --("11101111110000000000000000000000"),
         --("11101100100000001111110111101000"),
         --("10100010100000000000000000000110"),
         --("00000000000000000000000000000000"),
         --("01000000000000000000000000000000"),


         -- Filter sound test
         --("11101110100000000000000000100000"),
         --("11101110110000000000000100000000"),
         --("11101101100000000000111111111111"),
         --("00100111110000000000000000011001"),
         --("11101100100000001111001000110000"),
         --("10100010100000000000000000000101"),
         --("00000000000000000000000000000000"),
         --("11101101100000000000000000000000"),
         --("00100111110000000000000000011001"),
         --("11101100100000001111001000110000"),
         --("10100010100000000000000000001010"),
         --("00000000000000000000000000000000"),
         --("01000000000000000000000000000010"),

         -- Filter test sim
         --("11101110100000000000000010000010"),
         --("11101110110000000000000100000000"),
         --("11101101100000000010010100100101"),
         --("00000000000000000000000000000000"),
         --("00000000000000000000000000000000"),
         --("00000000000000000000000000000000"),
         --("00000000000000000000000000000000"),
         --("00000000000000000000000000000000"),
         --("11101101100000000010001100100011"),
         --("00000000000000000000000000000000"),
         --("00000000000000000000000000000000"),
         --("00000000000000000000000000000000"),
         --("00000000000000000000000000000000"),
         --("00000000000000000000000000000000"),
         --("11101101100000000010000000100000"),


         -- Test midi on/off
         --("11101000100000000000000000000000"),
         --("00100111110000000000000000000010"),
         --("11101100100000001111110111101000"),
         --("10100010100000000000000000000011"),
         --("00000000000000000000000000000000"),
         --("11101111110000000000000000000000"),
         --("11101100100000001111110111101000"),
         --("10100010100000000000000000000111"),
         --("00000000000000000000000000000000"),
         --("10100011100000000000000000000001"),
         --("00000000000000000000000000000000"),
         --("00100000010000000000000000011101"),
         --("00110010000000100000000000010000"),
         --("00110011010000100000000000010000"),
         --("10100000000000000000000000000000"),
         --("00000000000000000000000000000000"),
         --("11101000100000000000111111111111"),
         --("01000000000000000000000000000001"),
         --("00000000000000000000000000000000"),
      others =>
         ("00000" & "000" & "0000" & "0000" & "0000" & "0000" & "0000" & "0000")
      );
      
end pmemContent;
