package sout_constants is
   constant SOUT_CLK_FREQ  		: natural := 2268;
   constant SOUT_CLK_FREQ_WIDTH  : natural := 12; -- up to 4096
   constant SAMPLE_SIZE          : natural := 16;
   constant SAMPLE_SIZE_WIDTH    : natural := 6; 
end sout_constants;