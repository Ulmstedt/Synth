package MidiConstants is
    constant UART_CLK_PERIOD  : natural := 32;
    constant MIDI_WIDTH       : natural := 8;
end MidiConstants;