package MidiConstants is
    constant UART_CLK_PERIOD  : natural := 32;
    constant M1_WIDTH         : natural := 10;
    constant MIDI_WIDTH       : natural := 8;
end MidiConstants;