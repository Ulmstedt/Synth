package LCDConstants is

   constant XCOUNT_BITS          : natural =: 10;
   constant YCOUNT_BITS          : natural =: 9;

   constant tHA                  : natural =: 480;
   constant tHB                  : natural =: 45;
   
   constant tVA                  : natural =: 272;
   constant tVB                  : natural =: 16;

end LCDConstants;
