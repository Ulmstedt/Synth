library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

use work.records.all;


package pmemContent is
   constant pmemc : pmem_t := (
         ("00000" & "000" & "0000" & "0000" & "0000" & "0000" & "0000" & "0000"),
         ("11100" & "000" & "0000" & "0000" & "0000" & "0000" & "0000" & "0000"),
         ("00100" & "001" & "0000" & "0000" & "0000" & "0000" & "0000" & "0000"),
         ("01000" & "000" & "0000" & "0000" & "0000" & "0000" & "0000" & "0000"),
         ("00000" & "000" & "0000" & "0000" & "0000" & "0000" & "0000" & "0000"),
         ("00000" & "000" & "0000" & "0000" & "0000" & "0000" & "0000" & "0000"),
         ("00000" & "000" & "0000" & "0000" & "0000" & "0000" & "0000" & "0000"),
         ("01000" & "000" & "0000" & "0000" & "0000" & "0000" & "0000" & "0000"),
      others =>
         ("00000" & "000" & "0000" & "0000" & "0000" & "0000" & "0000" & "0000")
      );
      
end pmemContent;