package TouchConstants is
   constant VOLTAGE_WIDTH  : natural := 12;
   constant COORD_WIDTH    : natural := 9;
   constant MESSAGE_WIDTH  : natural := 15;
end TouchConstants;
