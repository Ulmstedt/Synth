library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

use work.records.all;


package pmemContent is

   constant pmemc : pmem_t := (
         ("11000" & "000" & "0000" & "0001" & "0000" & "0000" & "0000" & "0001"), -- STORE.c 1,#1
         ("11100" & "00001" & "000" & "0000" & "0000" & "000" & "0000" & "0001"), -- LOAD.a R1,1
         ("00110" & "00001" & "00001" & "0" & "0000" & "0000" & "0000" & "1000"), -- ADD R1,#8
         ("00100" & "00010" & "00" & "0000" & "0000" & "0000" & "000" & "00001"), -- MOVE R2,R1

         ("11001" & "000" & "0000" & "0010" & "0000" & "0000" & "000" & "00010"), -- STORE.r 2,R2
         ("00000" & "000" & "0000" & "0000" & "0000" & "0000" & "0000" & "0000"), -- NOP
         ("00000" & "000" & "0000" & "0000" & "0000" & "0000" & "0000" & "0000"), -- NOP
         ("11101" & "00001" & "000" & "0000" & "0000" & "000" & "0000" & "0100"), -- LOAD.c R1,4

         ("11101" & "00010" & "000" & "0000" & "0000" & "000" & "0000" & "1000"), -- LOAD.c R2,8
         ("00000" & "000" & "0000" & "0000" & "0000" & "0000" & "0000" & "0000"), -- NOP
         ("00000" & "000" & "0000" & "0000" & "0000" & "0000" & "0000" & "0000"), -- NOP
         ("00000" & "000" & "0000" & "0000" & "0000" & "0000" & "0000" & "0000"), -- NOP
         ("11010" & "000" & "0000" & "1000" & "000" & "0000" & "0001" & "00001"), -- STORE.wo 8,1,R1
         ("11011" & "000" & "0000" & "1000" & "00" & "0000" & "00001" & "00010"), -- STORE.wofr 8,R1,R2
         ("00000" & "000" & "0000" & "0000" & "0000" & "0000" & "0000" & "0000"), -- NOP

         --LOAD WITH OFFSET AND LOAD WITH OFFSET IN REGISTER LEFT TO TEST

      others =>
         ("00000" & "000" & "0000" & "0000" & "0000" & "0000" & "0000" & "0000")
      );
      
end pmemContent;
