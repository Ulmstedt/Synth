library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

use work.records.all;


package pmemContent is
   -- The content of the program memory
   constant pmemc : pmem_t := (
         ("11101100100000000000100000000000"),
         ("11101100110000001111110111101000"),
         ("11101000000000000000000000001010"),
         ("11101000100000000000000000001010"),
         ("00110001110000000000000000001000"),
         ("00110001110001000000000000001000"),
         ("11101000010000000000000000000000"),
         ("00101001010000000000000000000010"),
         ("00000000000000000000000000000000"),
         ("11011001111111110000000000000001"),
         ("00000000000000000000000000000000"),
         ("00110001000000000000000000000001"),
         ("00110011000000000000000000000000"),
         ("00000000000000000000000000000000"),
         ("10100000000000000000000000001000"),
         ("00000000000000000000000000000000"),
         ("11000001111101000000000110100101"),
         ("11000001111101010111111111111111"),
         ("10000011100000000000000000011010"),
         ("00000000000000000000000000000000"),
         ("10000010100000000000000010001011"),
         ("00000000000000000000000000000000"),
         ("10000011000000000000000010110110"),
         ("00000000000000000000000000000000"),
         ("01000000000000000000000000010010"),
         ("00000000000000000000000000000000"),
         ("00100010100000000000000000011101"),
         ("00110001100101000000000000001100"),
         ("00100000000000000000000000011101"),
         ("00110010000000000000000011111111"),
         ("00100000010000000000000000011110"),
         ("00110011000101000000000000001011"),
         ("10000000000000000000000001010001"),
         ("00000000000000000000000000000000"),
         ("00110011000101000000000000001110"),
         ("10000000000000000000000001100100"),
         ("00000000000000000000000000000000"),
         ("00110011000000000000000001010100"),
         ("10000000000000000000000010001000"),
         ("00000000000000000000000000000000"),
         ("11101001010000000000000000001010"),
         ("11101000100000000000001000000000"),
         ("00110011000000100000000000000000"),
         ("10000000000000000000000001000000"),
         ("00000000000000000000000000000000"),
         ("00110011000010100000000000000000"),
         ("10000000000000000000000001001111"),
         ("00000000000000000000000000000000"),
         ("11111001000001000000000000000000"),
         ("00110011000010000000000000000000"),
         ("10000000000000000000000000111000"),
         ("00000000000000000000000000000000"),
         ("00110000110010100000000000000001"),
         ("00110000010001000000000000001010"),
         ("01000000000000000000000000101101"),
         ("00000000000000000000000000000000"),
         ("11011000000000000001000000000000"),
         ("11101001000000000000000000000000"),
         ("11011000000000010001000000000100"),
         ("11101001000000000000100000000000"),
         ("11011000000000100001000000000100"),
         ("00110000100100000000000000000001"),
         ("01000000000000000000000001001111"),
         ("00000000000000000000000000000000"),
         ("00110011000010100000000000000000"),
         ("10000000000000000000000001001111"),
         ("00000000000000000000000000000000"),
         ("11111000110001000000000000000000"),
         ("00101011000000000000000000000011"),
         ("10100000000000000000000001001011"),
         ("00000000000000000000000000000000"),
         ("11101001000000000000000000000000"),
         ("00000000000000000000000000000000"),
         ("11011000000000000001000000000100"),
         ("00110001000100000000000000000001"),
         ("00110000110010100000000000000001"),
         ("00110000010001000000000000001010"),
         ("01000000000000000000000001000000"),
         ("00000000000000000000000000000000"),
         ("01000000000000000000000000010100"),
         ("00000000000000000000000000000000"),
         ("00110011000000000000000000000001"),
         ("10000000000000000000000001011001"),
         ("00000000000000000000000000000000"),
         ("00110011000000000000000000000111"),
         ("10000000000000000000000001011110"),
         ("00000000000000000000000000000000"),
         ("01000000000000000000000000010100"),
         ("00000000000000000000000000000000"),
         ("00100001000000000000000000000001"),
         ("00110001110010000000000000001000"),
         ("11001001111101000000000000000100"),
         ("01000000000000000000000000010100"),
         ("00000000000000000000000000000000"),
         ("11101001000000000000000001111111"),
         ("00101001000010000000000000000001"),
         ("00110001110010000000000000001000"),
         ("11001001111101010000000000000100"),
         ("01000000000000000000000000010100"),
         ("00000000000000000000000000000000"),
         ("00110011000101100000000000000000"),
         ("10000000000000000000000001101111"),
         ("00000000000000000000000000000000"),
         ("00110011000000100000000001111111"),
         ("10000000000000000000000001111101"),
         ("00000000000000000000000000000000"),
         ("00110011000000100000000000000000"),
         ("10000000000000000000000010000001"),
         ("00000000000000000000000000000000"),
         ("01000000000000000000000000010100"),
         ("00000000000000000000000000000000"),
         ("00110011000000100000000001111111"),
         ("10000000000000000000000001110111"),
         ("00000000000000000000000000000000"),
         ("00110011000000100000000000000000"),
         ("10000000000000000000000001111010"),
         ("00000000000000000000000000000000"),
         ("01000000000000000000000000010100"),
         ("00000000000000000000000000000000"),
         ("00110000101110000000000000000001"),
         ("01000000000000000000000000010100"),
         ("00000000000000000000000000000000"),
         ("00110001001110000000000000000001"),
         ("01000000000000000000000000010100"),
         ("00000000000000000000000000000000"),
         ("00110000100110000000000000000001"),
         ("00110010000110000000000000000011"),
         ("01000000000000000000000010000011"),
         ("00000000000000000000000000000000"),
         ("00110001000110000000000000000001"),
         ("00110010000110000000000000000011"),
         ("00100011010000000000000000001100"),
         ("00110001110110100000000000001000"),
         ("00110001010110100100000000000000"),
         ("01000000000000000000000000010100"),
         ("00000000000000000000000000000000"),
         ("00101010110101100000000000001011"),
         ("01000000000000000000000000010100"),
         ("00000000000000000000000000000000"),
         ("11101000100000000000001000000000"),
         ("11101001010000000000000000001010"),
         ("11101010010000000000000000000000"),
         ("11111000000001000000000000000000"),
         ("00110011000000000000000000000000"),
         ("10000000000000000000000010100101"),
         ("00000000000000000000000000000000"),
         ("11111001100000000000000000000000"),
         ("11111001110001000000000000000001"),
         ("00110000100011100000000000000001"),
         ("00101100010011000000000000000111"),
         ("00110011110011000000000000000110"),
         ("10000000000000000000000010011010"),
         ("00000000000000000000000000000000"),
         ("11101001110000000000000000000000"),
         ("00110000100001000000000000000001"),
         ("11011000000000000001000000000111"),
         ("00110001000001000000000000000001"),
         ("00110010000011000000000000111111"),
         ("00101000100011000000000000001101"),
         ("11111001000011000000000001010100"),
         ("00110011110010000000000000001111"),
         ("10000000000000000000000010100100"),
         ("00110001100010000000000000000100"),
         ("00110010010010001111000000000000"),
         ("00101000100100100000000000000100"),
         ("00110000100001000000000000001010"),
         ("00110001000010100000000000000001"),
         ("00110011000010100000000000000000"),
         ("10100000000000000000000010001110"),
         ("00000000000000000000000000000000"),
         ("11100110100000000000000111110100"),
         ("11100110110000000000000111110101"),
         ("00000000000000000000000000000000"),
         ("00000000000000000000000000000000"),
         ("00100101100000000000000000001001"),
         ("00000000000000000000000000000000"),
         ("00000000000000000000000000000000"),
         ("00000000000000000000000000000000"),
         ("00000000000000000000000000000000"),
         ("00100111110000000000000000011001"),
         ("01000000000000000000000000010110"),
         ("00000000000000000000000000000000"),
         ("11101100110000001111110111101000"),
         ("00110011000110000000000000000000"),
         ("10000000000000000000000011100111"),
         ("00000000000000000000000000000000"),
         ("00110011000110000000000000000001"),
         ("10000000000000000000000011101011"),
         ("00000000000000000000000000000000"),
         ("00110011000110000000000000000010"),
         ("10000000000000000000000011101111"),
         ("00000000000000000000000000000000"),
         ("00110011000110000000000000000011"),
         ("10000000000000000000000011110011"),
         ("00000000000000000000000000000000"),
         ("00100001000000000000000000011100"),
         ("00110010000010000000000000000011"),
         ("00110011000010000000000000000000"),
         ("10000000000000000000000011110111"),
         ("00000000000000000000000000000000"),
         ("00110011000010000000000000000001"),
         ("10000000000000000000000011111011"),
         ("00000000000000000000000000000000"),
         ("00110011000010000000000000000010"),
         ("10000000000000000000000011111111"),
         ("00000000000000000000000000000000"),
         ("00110011000010000000000000000011"),
         ("10000000000000000000000100000011"),
         ("00000000000000000000000000000000"),
         ("11100001000000000000000111110100"),
         ("00100001010000000000000000000100"),
         ("00110010000010001111000000000000"),
         ("00110001100010000000000000000100"),
         ("00100000000000000000000000000101"),
         ("00110001100000000000000000001000"),
         ("00110010000000000000000000001111"),
         ("00101000100010000000000000000000"),
         ("11001011010100000000000000000100"),
         ("11100001000000000000000111110101"),
         ("11101001010000000111111100000000"),
         ("00101001000010100000000000000100"),
         ("00100001000000000000000000000101"),
         ("00110010000010001111000000000000"),
         ("00110001100010000000000000000100"),
         ("00100000000000000000000000000101"),
         ("00110001100000000000000000001000"),
         ("00110010000000000000000000001111"),
         ("00101000100010000000000000000000"),
         ("11001011011011100000000000000100"),
         ("01000000000000000000000000011000"),
         ("00000000000000000000000000000000"),
         ("11000011000101000001100000010110"),
         ("11000011000101010001011100011110"),
         ("01000000000000000000000011000011"),
         ("00000000000000000000000000000000"),
         ("11000011000101000001100000010001"),
         ("11000011000101010001001100011110"),
         ("01000000000000000000000011000011"),
         ("00000000000000000000000000000000"),
         ("11000011000101000001100000001010"),
         ("11000011000101010001110000011110"),
         ("01000000000000000000000011000011"),
         ("00000000000000000000000000000000"),
         ("11000011000101000001100100010111"),
         ("11000011000101010001000100011110"),
         ("01000000000000000000000011000011"),
         ("00000000000000000000000000000000"),
         ("11000011001100100001001000010101"),
         ("11000011001100110001111000011110"),
         ("01000000000000000000000011010001"),
         ("00000000000000000000000000000000"),
         ("11000011001100100001000000010101"),
         ("11000011001100110001111000011110"),
         ("01000000000000000000000011010001"),
         ("00000000000000000000000000000000"),
         ("11000011001100100000101100010101"),
         ("11000011001100110001111000011110"),
         ("01000000000000000000000011010001"),
         ("00000000000000000000000000000000"),
         ("11000011001100100001001100010100"),
         ("11000011001100110001001100001110"),
         ("01000000000000000000000011010001"),
         ("00000000000000000000000000000000"),

      others =>
         ("00000" & "000" & "0000" & "0000" & "0000" & "0000" & "0000" & "0000")
      );
      
end pmemContent;
