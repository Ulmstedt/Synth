
package FilterConstants is
   constant AUDIO_WIDTH : natural := 16;
end FilterConstants;
