library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;


entity Touch is
   port(

      
      clk      : in std_logic;
      rst      : in std_logic;

   );
end Touch;


architecture Behavioural of Touch is
  
   
begin 
 
end Behavioural;
