library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

use work.records.all;


package pmemContent is

   constant pmemc : pmem_t := (
         --("11101" & "10010" & "000" & "0000" & "0000" & "000" & "0011" & "1111"), -- LOAD.c R18,15
            ("11101000100000000000000000000000"),
            ("00100111110000000000000000000010"),
            ("11101100100000001111110111101000"),
            ("10100010100000000000000000000011"),
            ("00000000000000000000000000000000"),
            ("11101111110000000000000000000000"),
            ("11101100100000001111110111101000"),
            ("10100010100000000000000000000111"),
            ("00000000000000000000000000000000"),
            ("10100011100000000000000000000001"),
            ("00000000000000000000000000000000"),
            ("00100000010000000000000000011101"),
            ("00110010000000100000000000010000"),
            ("00110011010000100000000000010000"),
            ("10100000000000000000000000000000"),
            ("00000000000000000000000000000000"),
            ("11101000100000000000111111111111"),
            ("00000000000000000000000000000000"),

      others =>
         ("00000" & "000" & "0000" & "0000" & "0000" & "0000" & "0000" & "0000")
      );
      
end pmemContent;
