package Constants is
    constant PMEM_WIDTH : natural := 32;
    constant ADDR_WIDTH : natural := 11;
    constant PMEM_HEIGHT : natural := 1024;
end Constants;
