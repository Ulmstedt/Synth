library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

use work.records.all;
use work.Constants.all;


package memContent is
   constant memc : mem_t := (
      -- Wavetables
      ("0001010111110010"), -- C4
      ("0001011101000000"), -- C#4
      ("0001100010100010"), -- D4
      ("0001101000011001"), -- D#4
      ("0001101110100111"), -- E4
      ("0001110101001010"), -- F4
      ("0001111100001010"), -- F#4
      ("0010000011100010"), -- G4
      ("0010001011010101"), -- G#4
      ("0010010011101000"), -- A4
      ("0010011100011010"), -- A#4
      ("0010100101101101"), -- B4
      
      -- 64 step square wave
      ("0000000000000000"), 
      ("0000000000000000"), 
      ("0000000000000000"), 
      ("0000000000000000"), 
      ("0000000000000000"), 
      ("0000000000000000"), 
      ("0000000000000000"), 
      ("0000000000000000"), 
      ("0000000000000000"), 
      ("0000000000000000"), 
      ("0000000000000000"), 
      ("0000000000000000"), 
      ("0000000000000000"), 
      ("0000000000000000"), 
      ("0000000000000000"), 
      ("0000000000000000"), 
      ("0000000000000000"), 
      ("0000000000000000"), 
      ("0000000000000000"), 
      ("0000000000000000"), 
      ("0000000000000000"), 
      ("0000000000000000"), 
      ("0000000000000000"), 
      ("0000000000000000"), 
      ("0000000000000000"), 
      ("0000000000000000"), 
      ("0000000000000000"), 
      ("0000000000000000"), 
      ("0000000000000000"), 
      ("0000000000000000"), 
      ("0000000000000000"), 
      ("0000000000000000"), 
      ("1111111111111111"), 
      ("1111111111111111"), 
      ("1111111111111111"), 
      ("1111111111111111"), 
      ("1111111111111111"), 
      ("1111111111111111"), 
      ("1111111111111111"), 
      ("1111111111111111"), 
      ("1111111111111111"), 
      ("1111111111111111"), 
      ("1111111111111111"), 
      ("1111111111111111"), 
      ("1111111111111111"), 
      ("1111111111111111"), 
      ("1111111111111111"), 
      ("1111111111111111"), 
      ("1111111111111111"), 
      ("1111111111111111"), 
      ("1111111111111111"), 
      ("1111111111111111"), 
      ("1111111111111111"), 
      ("1111111111111111"), 
      ("1111111111111111"), 
      ("1111111111111111"), 
      ("1111111111111111"), 
      ("1111111111111111"), 
      ("1111111111111111"), 
      ("1111111111111111"), 
      ("1111111111111111"), 
      ("1111111111111111"), 
      ("1111111111111111"), 
      ("1111111111111111"), 
      -- 64 step sine wave
      ("1000110010001011"), 
      ("1001100011111000"), 
      ("1010010100100111"), 
      ("1011000011111011"), 
      ("1011110001010101"), 
      ("1100011100011100"), 
      ("1101000100110010"), 
      ("1101101010000001"), 
      ("1110001011110001"), 
      ("1110101001101100"), 
      ("1111000011100001"), 
      ("1111011001000000"), 
      ("1111101001111100"), 
      ("1111110110001001"), 
      ("1111111101100001"), 
      ("1111111111111111"), 
      ("1111111101100001"), 
      ("1111110110001001"), 
      ("1111101001111100"), 
      ("1111011001000000"), 
      ("1111000011100001"), 
      ("1110101001101100"), 
      ("1110001011110001"), 
      ("1101101010000001"), 
      ("1101000100110010"), 
      ("1100011100011100"), 
      ("1011110001010101"), 
      ("1011000011111011"), 
      ("1010010100100111"), 
      ("1001100011111000"), 
      ("1000110010001011"), 
      ("0111111111111111"), 
      ("0111001101110011"), 
      ("0110011100000110"), 
      ("0101101011010111"), 
      ("0100111100000011"), 
      ("0100001110101001"), 
      ("0011100011100010"), 
      ("0010111011001100"), 
      ("0010010101111101"), 
      ("0001110100001101"), 
      ("0001010110010010"), 
      ("0000111100011101"), 
      ("0000100110111110"), 
      ("0000010110000010"), 
      ("0000001001110101"), 
      ("0000000010011101"), 
      ("0000000000000000"), 
      ("0000000010011101"), 
      ("0000001001110101"), 
      ("0000010110000010"), 
      ("0000100110111110"), 
      ("0000111100011101"), 
      ("0001010110010010"), 
      ("0001110100001101"), 
      ("0010010101111101"), 
      ("0010111011001100"), 
      ("0011100011100010"), 
      ("0100001110101001"), 
      ("0100111100000011"), 
      ("0101101011010111"), 
      ("0110011100000110"), 
      ("0111001101110011"), 
      ("0111111111111111"), 
      -- 64 step saw wave
      ("1111101111111111"), 
      ("1111011111111111"), 
      ("1111001111111111"), 
      ("1110111111111111"), 
      ("1110101111111111"), 
      ("1110011111111111"), 
      ("1110001111111111"), 
      ("1101111111111111"), 
      ("1101101111111111"), 
      ("1101011111111111"), 
      ("1101001111111111"), 
      ("1100111111111111"), 
      ("1100101111111111"), 
      ("1100011111111111"), 
      ("1100001111111111"), 
      ("1011111111111111"), 
      ("1011101111111111"), 
      ("1011011111111111"), 
      ("1011001111111111"), 
      ("1010111111111111"), 
      ("1010101111111111"), 
      ("1010011111111111"), 
      ("1010001111111111"), 
      ("1001111111111111"), 
      ("1001101111111111"), 
      ("1001011111111111"), 
      ("1001001111111111"), 
      ("1000111111111111"), 
      ("1000101111111111"), 
      ("1000011111111111"), 
      ("1000001111111111"), 
      ("0111111111111111"), 
      ("0111101111111111"), 
      ("0111011111111111"), 
      ("0111001111111111"), 
      ("0110111111111111"), 
      ("0110101111111111"), 
      ("0110011111111111"), 
      ("0110001111111111"), 
      ("0101111111111111"), 
      ("0101101111111111"), 
      ("0101011111111111"), 
      ("0101001111111111"), 
      ("0100111111111111"), 
      ("0100101111111111"), 
      ("0100011111111111"), 
      ("0100001111111111"), 
      ("0011111111111111"), 
      ("0011101111111111"), 
      ("0011011111111111"), 
      ("0011001111111111"), 
      ("0010111111111111"), 
      ("0010101111111111"), 
      ("0010011111111111"), 
      ("0010001111111111"), 
      ("0001111111111111"), 
      ("0001101111111111"), 
      ("0001011111111111"), 
      ("0001001111111111"), 
      ("0000111111111111"), 
      ("0000101111111111"), 
      ("0000011111111111"), 
      ("0000001111111111"), 
      ("0000000000000000"), 
      -- Cordic
      --TILE_MAP_OFFSET =>
      --   ("0000" & "0001" & "0000" & "0001" ),
      --TILE_MAP_OFFSET + 4 =>
      --   ("0000" & "0001" & "0000" & "0001" ),
      others =>
         ("0000" & "0000" & "0000" & "0000" )
      );
      
end memContent;
