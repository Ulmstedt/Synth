library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

use work.records.all;


package pmemContent is

   constant pmemc : pmem_t := (
        
         ("11101110100000000000000010000010"),
         ("11101110110000000000000100000000"),
         ("11101101100000000010010100100101"),
         ("00000000000000000000000000000000"),
         ("00000000000000000000000000000000"),
         ("00000000000000000000000000000000"),
         ("00000000000000000000000000000000"),
         ("00000000000000000000000000000000"),
         ("11101101100000000010001100100011"),
         ("00000000000000000000000000000000"),
         ("00000000000000000000000000000000"),
         ("00000000000000000000000000000000"),
         ("00000000000000000000000000000000"),
         ("00000000000000000000000000000000"),
         ("11101101100000000010000000100000"),


         -- Test midi on/off
         --("11101000100000000000000000000000"),
         --("00100111110000000000000000000010"),
         --("11101100100000001111110111101000"),
         --("10100010100000000000000000000011"),
         --("00000000000000000000000000000000"),
         --("11101111110000000000000000000000"),
         --("11101100100000001111110111101000"),
         --("10100010100000000000000000000111"),
         --("00000000000000000000000000000000"),
         --("10100011100000000000000000000001"),
         --("00000000000000000000000000000000"),
         --("00100000010000000000000000011101"),
         --("00110010000000100000000000010000"),
         --("00110011010000100000000000010000"),
         --("10100000000000000000000000000000"),
         --("00000000000000000000000000000000"),
         --("11101000100000000000111111111111"),
         --("01000000000000000000000000000001"),
         --("00000000000000000000000000000000"),
      others =>
         ("00000" & "000" & "0000" & "0000" & "0000" & "0000" & "0000" & "0000")
      );
      
end pmemContent;
