library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

use work.records.all;
use work.Constants.all;


package memContent is
   constant memc : mem_t := (
      -- Wavetables (calculated in advance as: freq * wavetable_length / sample rate
      ("0000000101011111"), -- "C0"
      ("0000000101110100"),
      ("0000000110001010"),
      ("0000000110100010"),
      ("0000000110111010"),
      ("0000000111010101"),
      ("0000000111110000"),
      ("0000001000001110"),
      ("0000001000101101"),
      ("0000001001001111"),
      ("0000001001110010"),
      ("0000001010010111"),
      ("0000001010111110"),
      ("0000001011101000"),
      ("0000001100010100"),
      ("0000001101000011"),
      ("0000001101110101"),
      ("0000001110101010"),
      ("0000001111100001"),
      ("0000010000011100"),
      ("0000010001011011"),
      ("0000010010011101"),
      ("0000010011100100"),
      ("0000010100101110"),
      ("0000010101111100"),
      ("0000010111010000"),
      ("0000011000101000"),
      ("0000011010000111"),
      ("0000011011101010"),
      ("0000011101010011"),
      ("0000011111000010"),
      ("0000100000111001"),
      ("0000100010110110"),
      ("0000100100111010"),
      ("0000100111000111"),
      ("0000101001011100"),
      ("0000101011111001"),
      ("0000101110100000"),
      ("0000110001010001"),
      ("0000110100001101"),
      ("0000110111010011"),
      ("0000111010100110"),
      ("0000111110000100"),
      ("0001000001110001"),
      ("0001000101101100"),
      ("0001001001110100"),
      ("0001001110001110"),
      ("0001010010110111"),
      ("0001010111110010"),
      ("0001011100111111"),
      ("0001100010100001"),
      ("0001101000011011"),
      ("0001101110100110"),
      ("0001110101001101"),
      ("0001111100001000"),
      ("0010000011100010"),
      ("0010001011011000"),
      ("0010010011101001"),
      ("0010011100011100"),
      ("0010100101101111"),
      ("0010101111100100"),
      ("0010111001111110"),
      ("0011000101000010"),
      ("0011010000110110"),
      ("0011011101001100"),
      ("0011101010011010"),
      ("0011111000010000"),
      ("0100000111000100"),
      ("0100010110110000"),
      ("0100100111010010"),
      ("0100111000111001"),
      ("0101001011011110"),
      ("0101011111000111"),
      ("0101110011111100"),
      ("0110001010000100"),
      ("0110100001101100"),
      ("0110111010011000"),
      ("0111010100110011"),
      ("0111110000100000"),
      ("1000001110001001"),
      ("1000101101011111"),
      ("1001001110100100"),
      ("1001110001110010"),
      ("1010010110111100"), -- "B6"
      
      -- 64 step square wave("0000000000000000"), 
      ("0000000000000000"), 
      ("0000000000000000"), 
      ("0000000000000000"), 
      ("0000000000000000"), 
      ("0000000000000000"), 
      ("0000000000000000"), 
      ("0000000000000000"), 
      ("0000000000000000"), 
      ("0000000000000000"), 
      ("0000000000000000"), 
      ("0000000000000000"), 
      ("0000000000000000"), 
      ("0000000000000000"), 
      ("0000000000000000"), 
      ("0000000000000000"), 
      ("0000000000000000"), 
      ("0000000000000000"), 
      ("0000000000000000"), 
      ("0000000000000000"), 
      ("0000000000000000"), 
      ("0000000000000000"), 
      ("0000000000000000"), 
      ("0000000000000000"), 
      ("0000000000000000"), 
      ("0000000000000000"), 
      ("0000000000000000"), 
      ("0000000000000000"), 
      ("0000000000000000"), 
      ("0000000000000000"), 
      ("0000000000000000"), 
      ("0000000000000000"), 
      ("1111111110000000"), 
      ("1111111110000000"), 
      ("1111111110000000"), 
      ("1111111110000000"), 
      ("1111111110000000"), 
      ("1111111110000000"), 
      ("1111111110000000"), 
      ("1111111110000000"), 
      ("1111111110000000"), 
      ("1111111110000000"), 
      ("1111111110000000"), 
      ("1111111110000000"), 
      ("1111111110000000"), 
      ("1111111110000000"), 
      ("1111111110000000"), 
      ("1111111110000000"), 
      ("1111111110000000"), 
      ("1111111110000000"), 
      ("1111111110000000"), 
      ("1111111110000000"), 
      ("1111111110000000"), 
      ("1111111110000000"), 
      ("1111111110000000"), 
      ("1111111110000000"), 
      ("1111111110000000"), 
      ("1111111110000000"), 
      ("1111111110000000"), 
      ("1111111110000000"), 
      ("1111111110000000"), 
      ("1111111110000000"), 
      ("1111111110000000"), 
      ("1111111110000000"), 
      -- 64 step sin wave("1000110001000101"), 
      ("1001100010101100"), 
      ("1010010011010101"), 
      ("1011000010100011"), 
      ("1011101111111000"), 
      ("1100011010111001"), 
      ("1101000011001011"), 
      ("1101101000010101"), 
      ("1110001010000000"), 
      ("1110100111111000"), 
      ("1111000001101010"), 
      ("1111010111000110"), 
      ("1111100111111111"), 
      ("1111110100001011"), 
      ("1111111011100010"), 
      ("1111111110000000"), 
      ("1111111011100010"), 
      ("1111110100001011"), 
      ("1111100111111111"), 
      ("1111010111000110"), 
      ("1111000001101010"), 
      ("1110100111111000"), 
      ("1110001010000000"), 
      ("1101101000010101"), 
      ("1101000011001011"), 
      ("1100011010111001"), 
      ("1011101111111000"), 
      ("1011000010100011"), 
      ("1010010011010101"), 
      ("1001100010101100"), 
      ("1000110001000101"), 
      ("0111111111000000"), 
      ("0111001100111010"), 
      ("0110011011010011"), 
      ("0101101010101010"), 
      ("0100111011011100"), 
      ("0100001110000111"), 
      ("0011100011000110"), 
      ("0010111010110100"), 
      ("0010010101101010"), 
      ("0001110011111111"), 
      ("0001010110000111"), 
      ("0000111100010101"), 
      ("0000100110111001"), 
      ("0000010110000000"), 
      ("0000001001110100"), 
      ("0000000010011101"), 
      ("0000000000000000"), 
      ("0000000010011101"), 
      ("0000001001110100"), 
      ("0000010110000000"), 
      ("0000100110111001"), 
      ("0000111100010101"), 
      ("0001010110000111"), 
      ("0001110011111111"), 
      ("0010010101101010"), 
      ("0010111010110100"), 
      ("0011100011000110"), 
      ("0100001110000111"), 
      ("0100111011011100"), 
      ("0101101010101010"), 
      ("0110011011010011"), 
      ("0111001100111010"), 
      ("0111111110111111"), 
      -- 64 step saw wave("1111101110000010"), 
      ("1111011110000100"), 
      ("1111001110000110"), 
      ("1110111110001000"), 
      ("1110101110001010"), 
      ("1110011110001100"), 
      ("1110001110001110"), 
      ("1101111110010000"), 
      ("1101101110010010"), 
      ("1101011110010100"), 
      ("1101001110010110"), 
      ("1100111110011000"), 
      ("1100101110011010"), 
      ("1100011110011100"), 
      ("1100001110011110"), 
      ("1011111110100000"), 
      ("1011101110100010"), 
      ("1011011110100100"), 
      ("1011001110100110"), 
      ("1010111110101000"), 
      ("1010101110101010"), 
      ("1010011110101100"), 
      ("1010001110101110"), 
      ("1001111110110000"), 
      ("1001101110110010"), 
      ("1001011110110100"), 
      ("1001001110110110"), 
      ("1000111110111000"), 
      ("1000101110111010"), 
      ("1000011110111100"), 
      ("1000001110111110"), 
      ("0111111111000000"), 
      ("0111101111000010"), 
      ("0111011111000100"), 
      ("0111001111000110"), 
      ("0110111111001000"), 
      ("0110101111001010"), 
      ("0110011111001100"), 
      ("0110001111001110"), 
      ("0101111111010000"), 
      ("0101101111010010"), 
      ("0101011111010100"), 
      ("0101001111010110"), 
      ("0100111111011000"), 
      ("0100101111011010"), 
      ("0100011111011100"), 
      ("0100001111011110"), 
      ("0011111111100000"), 
      ("0011101111100010"), 
      ("0011011111100100"), 
      ("0011001111100110"), 
      ("0010111111101000"), 
      ("0010101111101010"), 
      ("0010011111101100"), 
      ("0010001111101110"), 
      ("0001111111110000"), 
      ("0001101111110010"), 
      ("0001011111110100"), 
      ("0001001111110110"), 
      ("0000111111111000"), 
      ("0000101111111010"), 
      ("0000011111111100"), 
      ("0000001111111110"), 
      ("0000000000000000"), 
      -- Cordic
      --TILE_MAP_OFFSET =>
      --   ("0000" & "0001" & "0000" & "0001" ),
      --TILE_MAP_OFFSET + 4 =>
      --   ("0000" & "0001" & "0000" & "0001" ),
      others =>
         ("0000" & "0000" & "0000" & "0000" )
      );
      
end memContent;
