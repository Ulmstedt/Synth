
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

use work.constants.all;
use work.records.all;
use work.memContent.all;
use work.tilemapContent.all;

--Z4 now inside of memory
entity Memory is
   port(
      addr        : in std_logic_vector(ADDR_WIDTH - 1 downto 0);
      outputZ4    : out std_logic_vector(REG_WIDTH - 1 downto 0);
      doWrite     : in std_logic;
      newValue    : in std_logic_vector(REG_WIDTH - 1 downto 0);
      clk         : in std_logic;

      tmpOut      : out std_logic_vector(REG_WIDTH/2 - 1 downto 0);

      tileXcnt    : in std_logic_vector(HIGHER_BITS - 1 downto 0);
      tileYcnt    : in std_logic_vector(HIGHER_BITS - 1 downto 0);
      tileMapOut  : out std_logic_vector(TILE_MEM_ADRESS_BITS - 1 downto 0)
      
   );
end Memory;

architecture Behavioral of Memory is
   signal mem              : mem_t := memc;
   signal tilemap          : tilemap_t := tilemapc;
   signal rema             : std_logic_vector(5 downto 0);
   signal helpTileMem      : std_logic_vector(0 to REG_WIDTH - 1);
   signal maxXcnt          : std_logic_vector(HIGHER_BITS - 1 downto 0); -- Max 30
   signal maxYcnt          : std_logic_vector(HIGHER_BITS - 1 downto 0); -- Max 17
   signal isTilemap        : std_logic;
   
begin
   process(clk) is
   begin
      if rising_edge(clk) then
         if isTilemap = '0' then
            outputZ4 <= mem(to_integer(unsigned(addr) mod MEM_HEIGHT));
         elsif isTilemap = '1' then
            outputZ4 <= tilemap(to_integer((unsigned(addr) - TILE_MAP_OFFSET) mod TILE_MAP_HEIGHT));
         end if;
         if doWrite = '1' then
            if isTilemap = '0' then
               mem(to_integer(unsigned(addr)) mod MEM_HEIGHT) <= newValue;
            elsif isTilemap = '1' then
               tilemap(to_integer((unsigned(addr) - TILE_MAP_OFFSET) mod TILE_MAP_HEIGHT)) <= newValue;
            end if;
         end if;
      end if;
   end process;

   isTilemap <= '1' when to_integer(unsigned(addr) mod MEM_HEIGHT) >= TILE_MAP_OFFSET else
                '0';
   
   --varje slot i mem tar 2 tiles
   --en rad på skärmen = 30 tiles
   --en kolumn på skärmen = 17 tiles
   --Antar att tilemappen ligger kontinuerligt med tile 0 som första tilen dvs från offseten dvs tilemap[0][0] (första indexet motsvara raden, andra kolumn) i adress mem(TILE_MAP_OFFSET) och innehållet i bitarna 14 downto 10 i den. tile 60 (minns att det är räknat från 0 alltså i tilemap[1][0] osv
   --Antar att det gäller heltals division t e x 5/3 = 1, 5 rem 3 = 2
   -- XXXX XXXX XXXX XXXX

   maxXcnt <= tileXcnt when to_integer(unsigned(tileXcnt)) <= 29 else std_logic_vector(to_unsigned(29,HIGHER_BITS));
   maxYcnt <= tileYcnt when to_integer(unsigned(tileYcnt)) <= 16 else std_logic_vector(to_unsigned(16,HIGHER_BITS)); 
   rema <= std_logic_vector(to_unsigned(to_integer(unsigned(maxXcnt)) rem 2, 6));
   helpTileMem <= tilemap(to_integer(unsigned(maxYcnt)) * 15 + to_integer(unsigned(maxXcnt)) / 2);
   
   
   tileMapOut  <= helpTilemem(3 to 7) when rema = "000000" else
                  helpTilemem(11 to 15) when rema = "000001"  else
                  (others => '0');
   
   --tmpOut <= (others => '0');
   
end Behavioral;

