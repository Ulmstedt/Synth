library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

use work.records.all;


package pmemContent is

   constant pmemc : pmem_t := (
("11101100100000000000100000000000"),
("11101100110000001111110111101000"),
("11101000000000000000000000001010"),
("11101000100000000000000000001010"),
("00110001110000000000000000001000"),
("00110001110001000000000000001000"),
("11101000010000000000000000000000"),
("00101001010000000000000000000010"),
("00000000000000000000000000000000"),
("11011001111111110000000000000001"),
("00000000000000000000000000000000"),
("00110001000000000000000000000001"),
("00110011000000000000000000000000"),
("00000000000000000000000000000000"),
("10100000000000000000000000001000"),
("00000000000000000000000000000000"),
("11000001111101000000000110100101"),
("11000001111101010111111111111111"),
("10000011100000000000000000011010"),
("00000000000000000000000000000000"),
("10000010100000000000000010001001"),
("00000000000000000000000000000000"),
("10000011000000000000000010101110"),
("00000000000000000000000000000000"),
("01000000000000000000000000010010"),
("00000000000000000000000000000000"),
("00100010100000000000000000011101"),
("00110001100101000000000000001100"),
("00100000000000000000000000011101"),
("00110010000000000000000011111111"),
("00100000010000000000000000011110"),
("00110011000101000000000000001011"),
("10000000000000000000000001001111"),
("00000000000000000000000000000000"),
("00110011000101000000000000001110"),
("10000000000000000000000001100010"),
("00000000000000000000000000000000"),
("00110011000000000000000001010100"),
("10000000000000000000000010000110"),
("00000000000000000000000000000000"),
("11101001010000000000000000001010"),
("11101000100000000000001000000000"),
("00110011000000100000000000000000"),
("10000000000000000000000000111111"),
("00000000000000000000000000000000"),
("00110011000010100000000000000000"),
("10000000000000000000000001001101"),
("00000000000000000000000000000000"),
("11111001000001000000000000000000"),
("00110011000010000000000000000000"),
("10000000000000000000000000111000"),
("00000000000000000000000000000000"),
("00110000110010100000000000000001"),
("00110000010001000000000000001010"),
("01000000000000000000000000101101"),
("00000000000000000000000000000000"),
("11011000000000000001000000000000"),
("11101001000000000000000000000000"),
("11011000000000010001000000000100"),
("11101001000000000000100000000000"),
("11011000000000100001000000000100"),
("01000000000000000000000001001101"),
("00000000000000000000000000000000"),
("00110011000010100000000000000000"),
("10000000000000000000000001001101"),
("00000000000000000000000000000000"),
("11111000110001000000000000000000"),
("00101011000000000000000000000011"),
("10100000000000000000000001001001"),
("00000000000000000000000000000000"),
("11101001000000000000000000000000"),
("00000000000000000000000000000000"),
("11011000000000000001000000000100"),
("00110000110010100000000000000001"),
("00110000010001000000000000001010"),
("01000000000000000000000000111111"),
("00000000000000000000000000000000"),
("01000000000000000000000000010100"),
("00000000000000000000000000000000"),
("00110011000000000000000000000001"),
("10000000000000000000000001010111"),
("00000000000000000000000000000000"),
("00110011000000000000000000000111"),
("10000000000000000000000001011100"),
("00000000000000000000000000000000"),
("01000000000000000000000000010100"),
("00000000000000000000000000000000"),
("00100001000000000000000000000001"),
("00110001110010000000000000001000"),
("11001001111101000000000000000100"),
("01000000000000000000000000010100"),
("00000000000000000000000000000000"),
("11101001000000000000000001111111"),
("00110001000010000000000000000001"),
("00110001110010000000000000001000"),
("11001001111101010000000000000100"),
("01000000000000000000000000010100"),
("00000000000000000000000000000000"),
("00110011000101100000000000000000"),
("10000000000000000000000001101101"),
("00000000000000000000000000000000"),
("00110011000000100000000001111111"),
("10000000000000000000000001111011"),
("00000000000000000000000000000000"),
("00110011000000100000000000000000"),
("10000000000000000000000001111111"),
("00000000000000000000000000000000"),
("01000000000000000000000000010100"),
("00000000000000000000000000000000"),
("00110011000000100000000001111111"),
("10000000000000000000000001110101"),
("00000000000000000000000000000000"),
("00110011000000100000000000000000"),
("10000000000000000000000001111000"),
("00000000000000000000000000000000"),
("01000000000000000000000000010100"),
("00000000000000000000000000000000"),
("00110000101110000000000000000001"),
("01000000000000000000000000010100"),
("00000000000000000000000000000000"),
("00110001001110000000000000000001"),
("01000000000000000000000000010100"),
("00000000000000000000000000000000"),
("00110000100110000000000000000001"),
("00110010000110000000000000000011"),
("01000000000000000000000010000001"),
("00000000000000000000000000000000"),
("00110001000110000000000000000001"),
("00110010000110000000000000000011"),
("00100011010000000000000000001100"),
("00110001110110100000000000001000"),
("00110001010110100100000000000000"),
("01000000000000000000000000010100"),
("00000000000000000000000000000000"),
("00110010110101100000000000000000"),
("01000000000000000000000000010100"),
("00000000000000000000000000000000"),
("11101000100000000000001000000000"),
("11101001010000000000000000001010"),
("11101010010000000000000000000000"),
("11111000000001000000000000000000"),
("00110011000000000000000000000000"),
("10000000000000000000000010011101"),
("00000000000000000000000000000000"),
("11111001100000000000000000000000"),
("11111001110001000000000000000001"),
("00110000100011100000000000000001"),
("00101100010011000000000000000111"),
("00110000100001000000000000000001"),
("11011000000000000001000000000111"),
("00110001000001000000000000000001"),
("00110010000011000000000000111111"),
("00101000100011000000000000001101"),
("11111001000011000000000001010100"),
("11111000110001000000000000000010"),
("00101100010010000000000000000011"),
("00101000100100100000000000000100"),
("00110000100001000000000000001010"),
("00110001000010100000000000000001"),
("00110011000010100000000000000000"),
("10100000000000000000000010001100"),
("00000000000000000000000000000000"),
("11100110100000000000000111110100"),
("11100110110000000000000111110101"),
("00000000000000000000000000000000"),
("00000000000000000000000000000000"),
("00100101100000000000000000001001"),
("00000000000000000000000000000000"),
("00000000000000000000000000000000"),
("00000000000000000000000000000000"),
("00000000000000000000000000000000"),
("00100111110000000000000000011001"),
("01000000000000000000000000010110"),
("00000000000000000000000000000000"),
("11101100110000001111110111101000"),
("00110011000110000000000000000000"),
("10000000000000000000000011001011"),
("00000000000000000000000000000000"),
("00110011000110000000000000000001"),
("10000000000000000000000011001111"),
("00000000000000000000000000000000"),
("00110011000110000000000000000010"),
("10000000000000000000000011010011"),
("00000000000000000000000000000000"),
("00110011000110000000000000000011"),
("10000000000000000000000011010111"),
("00000000000000000000000000000000"),
("00100001000000000000000000011100"),
("00110010000010000000000000000011"),
("00110011000010000000000000000000"),
("10000000000000000000000011011011"),
("00000000000000000000000000000000"),
("00110011000010000000000000000001"),
("10000000000000000000000011011111"),
("00000000000000000000000000000000"),
("00110011000010000000000000000010"),
("10000000000000000000000011100011"),
("00000000000000000000000000000000"),
("00110011000010000000000000000011"),
("10000000000000000000000011100111"),
("00000000000000000000000000000000"),
("01000000000000000000000000011000"),
("00000000000000000000000000000000"),
("11001011001000100000000000010110"),
("11001011001000110000000000011110"),
("01000000000000000000000011001001"),
("00000000000000000000000000000000"),
("11001011001000100000000000010001"),
("11001011001000110000000000011110"),
("01000000000000000000000011001001"),
("00000000000000000000000000000000"),
("11001011001000100000000000001010"),
("11001011001000110000000000011110"),
("01000000000000000000000011001001"),
("00000000000000000000000000000000"),
("11001011001000100000000000010111"),
("11001011001000110000000000011110"),
("01000000000000000000000011001001"),
("00000000000000000000000000000000"),
("11001011010111100000000000010101"),
("11001011010111110000000000011110"),
("01000000000000000000000011001001"),
("00000000000000000000000000000000"),
("11001011010111100000000000010101"),
("11001011010111110000000000011110"),
("01000000000000000000000011001001"),
("00000000000000000000000000000000"),
("11001011010111100000000000010101"),
("11001011010111110000000000011110"),
("01000000000000000000000011001001"),
("00000000000000000000000000000000"),
("11001011010111100000000000010100"),
("11001011010111110000000000001110"),
("01000000000000000000000011001001"),
("00000000000000000000000000000000"),



         -- Simple sound test
         --("11101111110000000000111111111111"),
         --("11101100100000001111110111101000"),
         --("10100010100000000000000000000010"),
         --("00000000000000000000000000000000"),
         --("11101111110000000000000000000000"),
         --("11101100100000001111110111101000"),
         --("10100010100000000000000000000110"),
         --("00000000000000000000000000000000"),
         --("01000000000000000000000000000000"),


         -- Filter sound test
         --("11101110100000000000000000100000"),
         --("11101110110000000000000100000000"),
         --("11101101100000000000111111111111"),
         --("00100111110000000000000000011001"),
         --("11101100100000001111001000110000"),
         --("10100010100000000000000000000101"),
         --("00000000000000000000000000000000"),
         --("11101101100000000000000000000000"),
         --("00100111110000000000000000011001"),
         --("11101100100000001111001000110000"),
         --("10100010100000000000000000001010"),
         --("00000000000000000000000000000000"),
         --("01000000000000000000000000000010"),

         -- Filter test sim
         --("11101110100000000000000010000010"),
         --("11101110110000000000000100000000"),
         --("11101101100000000010010100100101"),
         --("00000000000000000000000000000000"),
         --("00000000000000000000000000000000"),
         --("00000000000000000000000000000000"),
         --("00000000000000000000000000000000"),
         --("00000000000000000000000000000000"),
         --("11101101100000000010001100100011"),
         --("00000000000000000000000000000000"),
         --("00000000000000000000000000000000"),
         --("00000000000000000000000000000000"),
         --("00000000000000000000000000000000"),
         --("00000000000000000000000000000000"),
         --("11101101100000000010000000100000"),


         -- Test midi on/off
         --("11101000100000000000000000000000"),
         --("00100111110000000000000000000010"),
         --("11101100100000001111110111101000"),
         --("10100010100000000000000000000011"),
         --("00000000000000000000000000000000"),
         --("11101111110000000000000000000000"),
         --("11101100100000001111110111101000"),
         --("10100010100000000000000000000111"),
         --("00000000000000000000000000000000"),
         --("10100011100000000000000000000001"),
         --("00000000000000000000000000000000"),
         --("00100000010000000000000000011101"),
         --("00110010000000100000000000010000"),
         --("00110011010000100000000000010000"),
         --("10100000000000000000000000000000"),
         --("00000000000000000000000000000000"),
         --("11101000100000000000111111111111"),
         --("01000000000000000000000000000001"),
         --("00000000000000000000000000000000"),
      others =>
         ("00000" & "000" & "0000" & "0000" & "0000" & "0000" & "0000" & "0000")
      );
      
end pmemContent;
