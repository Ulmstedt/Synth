library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

use work.records.all;


package pmemContent is

   constant pmemc : pmem_t := (
        
         ("11101110100000000000000010000010"),
         ("11101110110000000000000100000000"),
         ("11101101100000000010010100100101"),
         ("00000000000000000000000000000000"),
         ("00000000000000000000000000000000"),
         ("00000000000000000000000000000000"),
         ("00000000000000000000000000000000"),
         ("00000000000000000000000000000000"),
         ("11101101100000000010001100100011"),
         ("00000000000000000000000000000000"),
         ("00000000000000000000000000000000"),
         ("00000000000000000000000000000000"),
         ("00000000000000000000000000000000"),
         ("00000000000000000000000000000000"),
         ("11101101100000000010000000100000"),

      others =>
         ("00000" & "000" & "0000" & "0000" & "0000" & "0000" & "0000" & "0000")
      );
      
end pmemContent;
