library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

use work.records.all;


package pmemContent is

   constant pmemc : pmem_t := (
         --("11101" & "10010" & "000" & "0000" & "0000" & "000" & "0011" & "1111"), -- LOAD.c R18,15
            ("11101111110000001001001001001010"),
            ("11101100100000001100000011001110"),
            ("10100010100000000000000000000010"),
            ("00000000000000000000000000000000"),
            ("11101111110000001001001001001010"),
            ("11101100100000001100000011001110"),
            ("10100010100000000000000000000110"),
            ("00000000000000000000000000000000"),
            ("01000000000000000000000000000000"),

      others =>
         ("00000" & "000" & "0000" & "0000" & "0000" & "0000" & "0000" & "0000")
      );
      
end pmemContent;
