library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

use work.records.all;


package pmemContent is

   constant pmemc : pmem_t := (
         --program som räknar ut 0+1+2+3+4+5 = 15 och lägger resultatet i R2 
         ("11101" & "000" & "0000" & "0000" & "0000" & "0000" & "0000" & "0000"), -- LOAD.c R0,0
         ("11101" & "000" & "0100" & "0000" & "0000" & "0000" & "0000" & "0101"), -- LOAD.c R1,5
         ("00101" & "000" & "0100" & "0000" & "0000" & "0000" & "0000" & "0001"), -- ADDuns R0, R1
         ("00110" & "000" & "1100" & "0010" & "0000" & "0000" & "0000" & "0001"), -- SUBuns R1, 1
         ("00110" & "011" & "0000" & "0010" & "0000" & "0000" & "0000" & "0000"), -- CMP R1, 0
         ("10100" & "000" & "0000" & "0010" & "0000" & "0000" & "0000" & "0010"), -- BNCC(branch if Zero flag is not set) to $2
         ("00100" & "000" & "1000" & "0000" & "0000" & "0000" & "0000" & "0000"), -- MOVE R2,R0 
      others =>
         ("00000" & "000" & "0000" & "0000" & "0000" & "0000" & "0000" & "0000")
      );
      
end pmemContent;
