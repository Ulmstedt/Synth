library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

use work.records.all;


package pmemContent is

   constant pmemc : pmem_t := (
         ("11101" & "000" & "0100" & "0000" & "000" & "0000" & "0000" & "00100"), -- LOAD.c R1, 4
         ("00000" & "000" & "0000" & "0000" & "0000" & "0000" & "0000" & "0000"), --nop
         ("00000" & "000" & "0000" & "0000" & "0000" & "0000" & "0000" & "0000"),
         ("00000" & "000" & "0000" & "0000" & "0000" & "0000" & "0000" & "0000"),
         ("11010" & "000" & "0000" & "1000" & "000" & "0000" & "0001" & "00001"), -- ST.wo $8, 1,R1 
      others =>
         ("00000" & "000" & "0000" & "0000" & "0000" & "0000" & "0000" & "0000")
      );
      
end pmemContent;
